module test_master(a,b,c);
input a,b;
output c;

assign c =  a+b;

endmodule
